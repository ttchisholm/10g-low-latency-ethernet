package eg_frames;

logic [63:0] eg_tx_data[$] = {
64'h0707070707070707,
64'hd5555555555555fb,
64'h8b0e380577200008,
64'h0045000800000000,
64'h061b0000661c2800,
64'h00004d590000d79e,
64'h0000eb4a2839d168,
64'h12500c7a00007730,
64'h000000008462d21e,
64'h79f7eb9300000000,
64'h07070707070707fd,
64'h0707070707070707};

logic [7:0] eg_tx_ctl[$] = {
    8'b11111111,
    8'b00000001,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b00000000,
    8'b11111111,
    8'b11111111
};


logic [63:0] eg_rx_data[$] = {
    64'h000000000000001e,
    64'hd555555555555578,
    64'h8b0e380577200008,
    64'h0045000800000000,
    64'h061b0000661c2800,
    64'h00004d590000d79e,
    64'h0000eb4a2839d168,
    64'h12500c7a00007730,
    64'h000000008462d21e,
    64'h79f7eb9300000000,
    64'h0000000000000087
};

logic [1:0] eg_rx_header[$] = {
    2'b01,
    2'b01,
    2'b10,
    2'b10,
    2'b10,
    2'b10,
    2'b10,
    2'b10,
    2'b10,
    2'b10,
    2'b01
};

endpackage