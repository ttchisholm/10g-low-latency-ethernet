package eg_frames;

logic [31:0] eg_tx_data[$] = {
32'h07070707,
32'h07070707,
32'hfb555555,
32'h555555d5,
32'h08002077,
32'h05380e8b,
32'h00000000,
32'h08004500,
32'h00281c66,
32'h00001b06,
32'h9ed70000,
32'h594d0000,
32'h68d13928,
32'h4aeb0000,
32'h30770000,
32'h7a0c5012,
32'h1ed26284,
32'h00000000,
32'h00000000,
32'h93ebf779,
32'hfd070707,
32'h07070707};

logic [3:0] eg_tx_ctl[$] = {
    4'b1111,
    4'b1111,
    4'b1000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b0000,
    4'b1111,
    4'b1111
};

endpackage